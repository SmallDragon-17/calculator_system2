module MULTI2TEST;


  reg [1:0] a;
  reg [1:0] b;
  wire [3:0] s;
  integer i, j, k, m;
  //reg a1,a0,b1,b0;
  //wire d3,d2,d1,d0;

  MULTI2 bbb(a,b,s);
    initial begin
      $dumpfile("mulit2test.vcd");
      $dumpvars(0,MULTI2TEST);
      $monitor("%t: a1 = %b, a0 = %b,b1 = %b, b0 = %b, d3 = %b, d2 = %b, d1 = %b, d0 = %b", $time, a[1],a[0],b[1],b[0],s[3],s[2],s[1],s[0]);

       a[1]=0; a[0]=0; b[1]=0; b[0]=0;
      // a = 2'b00; b = 2'b00;
      // b[1] = 0; b[0] = 0;
      // for (i = 0; i < 2; i = i + 1)
      //   for (k = 0; k < 2; k = k + 1)
      //     for (m = 0; m < 2; m = m + 1) begin
      //       #10 b[0] = i; a[1] = k; a[0] = m;
      //     end
      for(i=0; i<2; i=i+1) 
        for(j=0; j<2; j=j+1)
          for(k=0; k<2; k=k+1)
            for(m=0; m<2; m=m+1) begin
              #10 b[0] = j; b[1] = i; a[0] = m; a[1] = k;
            end

      //   a[1]=0; a[0]=0; b[1]=0; b[0]=0;
      // #10 a[1]=0; a[0]=1; b[1]=0; b[0]=0;
      // #10 a[1]=1; a[0]=0; b[1]=0; b[0]=0;
      // #10 a[1]=1; a[0]=1; b[1]=0; b[0]=0;
      // #10 a[1]=0; a[0]=0; b[1]=0; b[0]=1;
      // #10 a[1]=0; a[0]=1; b[1]=0; b[0]=1;
      // #10 a[1]=1; a[0]=0; b[1]=0; b[0]=1;
      // #10 a[1]=1; a[0]=1; b[1]=0; b[0]=1;
      // #10 a[1]=0; a[0]=0; b[1]=1; b[0]=0;
      // #10 a[1]=0; a[0]=1; b[1]=1; b[0]=0;
      // #10 a[1]=1; a[0]=0; b[1]=1; b[0]=0;
      // #10 a[1]=1; a[0]=1; b[1]=1; b[0]=0;
      // #10 a[1]=0; a[0]=0; b[1]=1; b[0]=1;
      // #10 a[1]=0; a[0]=1; b[1]=1; b[0]=1;
      // #10 a[1]=1; a[0]=0; b[1]=1; b[0]=1;
      // #10 a[1]=1; a[0]=1; b[1]=1; b[0]=1;
      #10 $finish;
    end
endmodule 

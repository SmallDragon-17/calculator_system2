module OR2(A,B,X);

input A,B;
output X;

assign X = A | B;

endmodule

